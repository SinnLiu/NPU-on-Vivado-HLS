module pe_acc(
    input  [1023:0] mult_result,
    output [31:0]   acc_result
  );
  genvar i;
  genvar j;
  wire [31:0] int16_result[31:0][5:0];
  /* add tree */
  // TODO:
endmodule
